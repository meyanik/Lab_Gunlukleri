magic
tech sky130A
magscale 1 2
timestamp 1658993734
<< nwell >>
rect -596 -2573 596 2573
<< pmoslvt >>
rect -400 1354 400 2354
rect -400 118 400 1118
rect -400 -1118 400 -118
rect -400 -2354 400 -1354
<< pdiff >>
rect -458 2342 -400 2354
rect -458 1366 -446 2342
rect -412 1366 -400 2342
rect -458 1354 -400 1366
rect 400 2342 458 2354
rect 400 1366 412 2342
rect 446 1366 458 2342
rect 400 1354 458 1366
rect -458 1106 -400 1118
rect -458 130 -446 1106
rect -412 130 -400 1106
rect -458 118 -400 130
rect 400 1106 458 1118
rect 400 130 412 1106
rect 446 130 458 1106
rect 400 118 458 130
rect -458 -130 -400 -118
rect -458 -1106 -446 -130
rect -412 -1106 -400 -130
rect -458 -1118 -400 -1106
rect 400 -130 458 -118
rect 400 -1106 412 -130
rect 446 -1106 458 -130
rect 400 -1118 458 -1106
rect -458 -1366 -400 -1354
rect -458 -2342 -446 -1366
rect -412 -2342 -400 -1366
rect -458 -2354 -400 -2342
rect 400 -1366 458 -1354
rect 400 -2342 412 -1366
rect 446 -2342 458 -1366
rect 400 -2354 458 -2342
<< pdiffc >>
rect -446 1366 -412 2342
rect 412 1366 446 2342
rect -446 130 -412 1106
rect 412 130 446 1106
rect -446 -1106 -412 -130
rect 412 -1106 446 -130
rect -446 -2342 -412 -1366
rect 412 -2342 446 -1366
<< nsubdiff >>
rect -560 2503 -464 2537
rect 464 2503 560 2537
rect -560 2441 -526 2503
rect 526 2441 560 2503
rect -560 -2503 -526 -2441
rect 526 -2503 560 -2441
rect -560 -2537 -464 -2503
rect 464 -2537 560 -2503
<< nsubdiffcont >>
rect -464 2503 464 2537
rect -560 -2441 -526 2441
rect 526 -2441 560 2441
rect -464 -2537 464 -2503
<< poly >>
rect -400 2435 400 2451
rect -400 2401 -384 2435
rect 384 2401 400 2435
rect -400 2354 400 2401
rect -400 1307 400 1354
rect -400 1273 -384 1307
rect 384 1273 400 1307
rect -400 1257 400 1273
rect -400 1199 400 1215
rect -400 1165 -384 1199
rect 384 1165 400 1199
rect -400 1118 400 1165
rect -400 71 400 118
rect -400 37 -384 71
rect 384 37 400 71
rect -400 21 400 37
rect -400 -37 400 -21
rect -400 -71 -384 -37
rect 384 -71 400 -37
rect -400 -118 400 -71
rect -400 -1165 400 -1118
rect -400 -1199 -384 -1165
rect 384 -1199 400 -1165
rect -400 -1215 400 -1199
rect -400 -1273 400 -1257
rect -400 -1307 -384 -1273
rect 384 -1307 400 -1273
rect -400 -1354 400 -1307
rect -400 -2401 400 -2354
rect -400 -2435 -384 -2401
rect 384 -2435 400 -2401
rect -400 -2451 400 -2435
<< polycont >>
rect -384 2401 384 2435
rect -384 1273 384 1307
rect -384 1165 384 1199
rect -384 37 384 71
rect -384 -71 384 -37
rect -384 -1199 384 -1165
rect -384 -1307 384 -1273
rect -384 -2435 384 -2401
<< locali >>
rect -560 2503 -464 2537
rect 464 2503 560 2537
rect -560 2441 -526 2503
rect 526 2441 560 2503
rect -400 2401 -384 2435
rect 384 2401 400 2435
rect -446 2342 -412 2358
rect -446 1350 -412 1366
rect 412 2342 446 2358
rect 412 1350 446 1366
rect -400 1273 -384 1307
rect 384 1273 400 1307
rect -400 1165 -384 1199
rect 384 1165 400 1199
rect -446 1106 -412 1122
rect -446 114 -412 130
rect 412 1106 446 1122
rect 412 114 446 130
rect -400 37 -384 71
rect 384 37 400 71
rect -400 -71 -384 -37
rect 384 -71 400 -37
rect -446 -130 -412 -114
rect -446 -1122 -412 -1106
rect 412 -130 446 -114
rect 412 -1122 446 -1106
rect -400 -1199 -384 -1165
rect 384 -1199 400 -1165
rect -400 -1307 -384 -1273
rect 384 -1307 400 -1273
rect -446 -1366 -412 -1350
rect -446 -2358 -412 -2342
rect 412 -1366 446 -1350
rect 412 -2358 446 -2342
rect -400 -2435 -384 -2401
rect 384 -2435 400 -2401
rect -560 -2503 -526 -2441
rect 526 -2503 560 -2441
rect -560 -2537 -464 -2503
rect 464 -2537 560 -2503
<< viali >>
rect -384 2401 384 2435
rect -446 1366 -412 2342
rect 412 1366 446 2342
rect -384 1273 384 1307
rect -384 1165 384 1199
rect -446 130 -412 1106
rect 412 130 446 1106
rect -384 37 384 71
rect -384 -71 384 -37
rect -446 -1106 -412 -130
rect 412 -1106 446 -130
rect -384 -1199 384 -1165
rect -384 -1307 384 -1273
rect -446 -2342 -412 -1366
rect 412 -2342 446 -1366
rect -384 -2435 384 -2401
<< metal1 >>
rect -396 2435 396 2441
rect -396 2401 -384 2435
rect 384 2401 396 2435
rect -396 2395 396 2401
rect -452 2342 -406 2354
rect -452 1366 -446 2342
rect -412 1366 -406 2342
rect -452 1354 -406 1366
rect 406 2342 452 2354
rect 406 1366 412 2342
rect 446 1366 452 2342
rect 406 1354 452 1366
rect -396 1307 396 1313
rect -396 1273 -384 1307
rect 384 1273 396 1307
rect -396 1267 396 1273
rect -396 1199 396 1205
rect -396 1165 -384 1199
rect 384 1165 396 1199
rect -396 1159 396 1165
rect -452 1106 -406 1118
rect -452 130 -446 1106
rect -412 130 -406 1106
rect -452 118 -406 130
rect 406 1106 452 1118
rect 406 130 412 1106
rect 446 130 452 1106
rect 406 118 452 130
rect -396 71 396 77
rect -396 37 -384 71
rect 384 37 396 71
rect -396 31 396 37
rect -396 -37 396 -31
rect -396 -71 -384 -37
rect 384 -71 396 -37
rect -396 -77 396 -71
rect -452 -130 -406 -118
rect -452 -1106 -446 -130
rect -412 -1106 -406 -130
rect -452 -1118 -406 -1106
rect 406 -130 452 -118
rect 406 -1106 412 -130
rect 446 -1106 452 -130
rect 406 -1118 452 -1106
rect -396 -1165 396 -1159
rect -396 -1199 -384 -1165
rect 384 -1199 396 -1165
rect -396 -1205 396 -1199
rect -396 -1273 396 -1267
rect -396 -1307 -384 -1273
rect 384 -1307 396 -1273
rect -396 -1313 396 -1307
rect -452 -1366 -406 -1354
rect -452 -2342 -446 -1366
rect -412 -2342 -406 -1366
rect -452 -2354 -406 -2342
rect 406 -1366 452 -1354
rect 406 -2342 412 -1366
rect 446 -2342 452 -1366
rect 406 -2354 452 -2342
rect -396 -2401 396 -2395
rect -396 -2435 -384 -2401
rect 384 -2435 396 -2401
rect -396 -2441 396 -2435
<< properties >>
string FIXED_BBOX -543 -2520 543 2520
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 5.0 l 4.0 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
