magic
tech sky130A
magscale 1 2
timestamp 1659002813
<< nwell >>
rect 792 492 1214 1566
rect 1471 503 1893 1577
<< pwell >>
rect 808 146 1230 410
rect 680 61 1230 146
rect 737 -252 765 61
rect 808 -24 1230 61
rect 1515 62 1937 410
rect 2020 62 2121 391
rect 1515 27 2121 62
rect 808 -75 1259 -24
rect 1515 -37 1937 27
rect 1465 -63 1937 -37
rect 808 -210 1230 -75
rect 1500 -84 1937 -63
rect 1515 -210 1937 -84
rect 737 -314 1106 -252
rect 2020 -383 2121 27
rect 1281 -434 2146 -383
rect 1281 -436 1951 -434
rect 2020 -436 2121 -434
<< nmos >>
rect 1004 0 1034 200
rect 1711 0 1741 200
<< pmos >>
rect 988 1147 1018 1347
rect 988 711 1018 911
rect 1667 1158 1697 1358
rect 1667 722 1697 922
<< ndiff >>
rect 946 188 1004 200
rect 946 12 958 188
rect 992 12 1004 188
rect 946 0 1004 12
rect 1034 188 1092 200
rect 1034 12 1046 188
rect 1080 12 1092 188
rect 1034 0 1092 12
rect 1653 188 1711 200
rect 1653 12 1665 188
rect 1699 12 1711 188
rect 1653 0 1711 12
rect 1741 188 1799 200
rect 1741 12 1753 188
rect 1787 12 1799 188
rect 1741 0 1799 12
<< pdiff >>
rect 930 1335 988 1347
rect 930 1159 942 1335
rect 976 1159 988 1335
rect 930 1147 988 1159
rect 1018 1335 1076 1347
rect 1018 1159 1030 1335
rect 1064 1159 1076 1335
rect 1018 1147 1076 1159
rect 930 899 988 911
rect 930 723 942 899
rect 976 723 988 899
rect 930 711 988 723
rect 1018 899 1076 911
rect 1018 723 1030 899
rect 1064 723 1076 899
rect 1018 711 1076 723
rect 1609 1346 1667 1358
rect 1609 1170 1621 1346
rect 1655 1170 1667 1346
rect 1609 1158 1667 1170
rect 1697 1346 1755 1358
rect 1697 1170 1709 1346
rect 1743 1170 1755 1346
rect 1697 1158 1755 1170
rect 1609 910 1667 922
rect 1609 734 1621 910
rect 1655 734 1667 910
rect 1609 722 1667 734
rect 1697 910 1755 922
rect 1697 734 1709 910
rect 1743 734 1755 910
rect 1697 722 1755 734
<< ndiffc >>
rect 958 12 992 188
rect 1046 12 1080 188
rect 1665 12 1699 188
rect 1753 12 1787 188
<< pdiffc >>
rect 942 1159 976 1335
rect 1030 1159 1064 1335
rect 942 723 976 899
rect 1030 723 1064 899
rect 1621 1170 1655 1346
rect 1709 1170 1743 1346
rect 1621 734 1655 910
rect 1709 734 1743 910
<< psubdiff >>
rect 844 340 940 374
rect 1098 340 1194 374
rect 844 278 878 340
rect 1160 278 1194 340
rect 844 -140 878 -78
rect 1160 -140 1194 -78
rect 844 -174 940 -140
rect 1098 -174 1194 -140
rect 1551 340 1647 374
rect 1805 340 1901 374
rect 1551 278 1585 340
rect 1867 278 1901 340
rect 1551 -140 1585 -78
rect 1867 -140 1901 -78
rect 1551 -174 1647 -140
rect 1805 -174 1901 -140
<< nsubdiff >>
rect 828 1496 924 1530
rect 1082 1496 1178 1530
rect 828 1434 862 1496
rect 1144 1434 1178 1496
rect 828 562 862 624
rect 1144 562 1178 624
rect 828 528 924 562
rect 1082 528 1178 562
rect 1507 1507 1603 1541
rect 1761 1507 1857 1541
rect 1507 1445 1541 1507
rect 1823 1445 1857 1507
rect 1507 573 1541 635
rect 1823 573 1857 635
rect 1507 539 1603 573
rect 1761 539 1857 573
<< psubdiffcont >>
rect 940 340 1098 374
rect 844 -78 878 278
rect 1160 -78 1194 278
rect 940 -174 1098 -140
rect 1647 340 1805 374
rect 1551 -78 1585 278
rect 1867 -78 1901 278
rect 1647 -174 1805 -140
<< nsubdiffcont >>
rect 924 1496 1082 1530
rect 828 624 862 1434
rect 1144 624 1178 1434
rect 924 528 1082 562
rect 1603 1507 1761 1541
rect 1507 635 1541 1445
rect 1823 635 1857 1445
rect 1603 539 1761 573
<< poly >>
rect 970 1428 1036 1444
rect 970 1394 986 1428
rect 1020 1394 1036 1428
rect 970 1378 1036 1394
rect 988 1347 1018 1378
rect 988 1116 1018 1147
rect 970 1100 1036 1116
rect 970 1066 986 1100
rect 1020 1066 1036 1100
rect 970 1050 1036 1066
rect 970 992 1036 1008
rect 970 958 986 992
rect 1020 958 1036 992
rect 970 942 1036 958
rect 988 911 1018 942
rect 988 680 1018 711
rect 970 664 1036 680
rect 970 630 986 664
rect 1020 630 1036 664
rect 970 614 1036 630
rect 1649 1439 1715 1455
rect 1649 1405 1665 1439
rect 1699 1405 1715 1439
rect 1649 1389 1715 1405
rect 1667 1358 1697 1389
rect 1667 1127 1697 1158
rect 1649 1111 1715 1127
rect 1649 1077 1665 1111
rect 1699 1077 1715 1111
rect 1649 1061 1715 1077
rect 1649 1003 1715 1019
rect 1649 969 1665 1003
rect 1699 969 1715 1003
rect 1649 953 1715 969
rect 1667 922 1697 953
rect 1667 691 1697 722
rect 1649 675 1715 691
rect 1649 641 1665 675
rect 1699 641 1715 675
rect 1649 625 1715 641
rect 986 272 1052 288
rect 986 238 1002 272
rect 1036 238 1052 272
rect 986 222 1052 238
rect 1004 200 1034 222
rect 1004 -22 1034 0
rect 986 -38 1052 -22
rect 986 -72 1002 -38
rect 1036 -72 1052 -38
rect 986 -88 1052 -72
rect 1693 272 1759 288
rect 1693 238 1709 272
rect 1743 238 1759 272
rect 1693 222 1759 238
rect 1711 200 1741 222
rect 1711 -22 1741 0
rect 1693 -38 1759 -22
rect 1693 -72 1709 -38
rect 1743 -72 1759 -38
rect 1693 -88 1759 -72
<< polycont >>
rect 986 1394 1020 1428
rect 986 1066 1020 1100
rect 986 958 1020 992
rect 986 630 1020 664
rect 1665 1405 1699 1439
rect 1665 1077 1699 1111
rect 1665 969 1699 1003
rect 1665 641 1699 675
rect 1002 238 1036 272
rect 1002 -72 1036 -38
rect 1709 238 1743 272
rect 1709 -72 1743 -38
<< locali >>
rect 828 1496 924 1530
rect 1082 1496 1178 1530
rect 828 1434 862 1496
rect 1144 1434 1178 1496
rect 970 1394 986 1428
rect 1020 1394 1036 1428
rect 942 1335 976 1351
rect 942 1143 976 1159
rect 1030 1335 1064 1351
rect 1030 1143 1064 1159
rect 970 1066 986 1100
rect 1020 1066 1036 1100
rect 970 958 986 992
rect 1020 958 1036 992
rect 942 899 976 915
rect 942 707 976 723
rect 1030 899 1064 915
rect 1030 707 1064 723
rect 970 630 986 664
rect 1020 630 1036 664
rect 828 562 862 624
rect 1144 562 1178 624
rect 828 528 924 562
rect 1082 528 1178 562
rect 1507 1507 1603 1541
rect 1761 1507 1857 1541
rect 1507 1445 1541 1507
rect 1823 1445 1857 1507
rect 1649 1405 1665 1439
rect 1699 1405 1715 1439
rect 1621 1346 1655 1362
rect 1621 1154 1655 1170
rect 1709 1346 1743 1362
rect 1709 1154 1743 1170
rect 1649 1077 1665 1111
rect 1699 1077 1715 1111
rect 1649 969 1665 1003
rect 1699 969 1715 1003
rect 1621 910 1655 926
rect 1621 718 1655 734
rect 1709 910 1743 926
rect 1709 718 1743 734
rect 1649 641 1665 675
rect 1699 641 1715 675
rect 1507 573 1541 635
rect 1823 573 1857 635
rect 1507 539 1603 573
rect 1761 539 1857 573
rect 844 340 940 374
rect 1098 340 1194 374
rect 844 278 878 340
rect 1160 280 1194 340
rect 1551 340 1647 374
rect 1805 340 1901 374
rect 986 238 1002 272
rect 1036 238 1052 272
rect 958 188 992 204
rect 958 -4 992 12
rect 1046 188 1080 204
rect 1046 -4 1080 12
rect 1551 278 1585 340
rect 1867 278 1901 340
rect 1693 238 1709 272
rect 1743 238 1759 272
rect 986 -72 1002 -38
rect 1036 -72 1052 -38
rect 844 -140 878 -78
rect 1160 -140 1194 -78
rect 844 -174 940 -140
rect 1098 -174 1194 -140
rect 1665 188 1699 204
rect 1665 -4 1699 12
rect 1753 188 1787 204
rect 1753 -4 1787 12
rect 1693 -72 1709 -38
rect 1743 -72 1759 -38
rect 1551 -140 1585 -78
rect 1867 -140 1901 -78
rect 1551 -174 1647 -140
rect 1805 -174 1901 -140
<< viali >>
rect 986 1394 1020 1428
rect 826 951 828 1191
rect 828 951 862 1191
rect 862 951 864 1191
rect 942 1159 976 1335
rect 1030 1159 1064 1335
rect 1143 1118 1144 1321
rect 1144 1118 1177 1321
rect 986 1066 1020 1100
rect 986 958 1020 992
rect 942 723 976 899
rect 1030 723 1064 899
rect 986 630 1020 664
rect 1665 1405 1699 1439
rect 1507 1124 1541 1327
rect 1621 1170 1655 1346
rect 1709 1170 1743 1346
rect 1665 1077 1699 1111
rect 1665 969 1699 1003
rect 1621 734 1655 910
rect 1709 734 1743 910
rect 1665 641 1699 675
rect 1160 278 1195 280
rect 845 -78 878 264
rect 878 -78 879 264
rect 1002 238 1036 272
rect 958 12 992 188
rect 1046 12 1080 188
rect 1160 132 1194 278
rect 1194 132 1195 278
rect 1551 195 1585 277
rect 1709 238 1743 272
rect 1002 -72 1036 -38
rect 1665 12 1699 188
rect 1753 12 1787 188
rect 1709 -72 1743 -38
<< metal1 >>
rect 680 1747 1393 1749
rect 680 1746 1436 1747
rect 680 1693 1397 1746
rect 1450 1693 1460 1746
rect 681 1691 1436 1693
rect 404 1111 604 1223
rect 681 1111 746 1691
rect 1217 1575 1227 1628
rect 1280 1627 1290 1628
rect 1280 1626 1698 1627
rect 2066 1626 2096 1628
rect 1280 1575 2096 1626
rect 1677 1574 2096 1575
rect 966 1439 1714 1460
rect 966 1428 1665 1439
rect 966 1394 986 1428
rect 1020 1405 1665 1428
rect 1699 1405 1714 1439
rect 1020 1394 1714 1405
rect 966 1389 1714 1394
rect 974 1388 1032 1389
rect 936 1335 982 1347
rect 820 1191 870 1203
rect 936 1196 942 1335
rect 904 1193 942 1196
rect 820 1112 826 1191
rect 790 1111 826 1112
rect 404 1051 826 1111
rect 404 1023 604 1051
rect 790 1049 826 1051
rect 820 951 826 1049
rect 864 1112 870 1191
rect 903 1159 942 1193
rect 976 1159 982 1335
rect 903 1147 982 1159
rect 1024 1335 1070 1347
rect 1615 1346 1661 1358
rect 1024 1159 1030 1335
rect 1064 1239 1070 1335
rect 1137 1321 1183 1333
rect 1064 1213 1095 1239
rect 1064 1159 1105 1213
rect 1024 1147 1105 1159
rect 903 1112 938 1147
rect 1058 1145 1105 1147
rect 864 1049 938 1112
rect 864 951 870 1049
rect 820 939 870 951
rect 903 911 938 1049
rect 970 1100 1034 1110
rect 970 1066 986 1100
rect 1020 1066 1034 1100
rect 970 992 1034 1066
rect 970 958 986 992
rect 1020 958 1034 992
rect 970 940 1034 958
rect 1074 1029 1105 1145
rect 1137 1118 1143 1321
rect 1177 1215 1183 1321
rect 1501 1327 1547 1339
rect 1501 1215 1507 1327
rect 1177 1181 1507 1215
rect 1177 1118 1183 1181
rect 1137 1106 1183 1118
rect 1501 1124 1507 1181
rect 1541 1124 1547 1327
rect 1615 1229 1621 1346
rect 1584 1218 1621 1229
rect 1583 1170 1621 1218
rect 1655 1170 1661 1346
rect 1583 1158 1661 1170
rect 1703 1346 1749 1358
rect 1703 1170 1709 1346
rect 1743 1298 1749 1346
rect 2066 1298 2096 1574
rect 1743 1205 2096 1298
rect 1743 1170 1749 1205
rect 1703 1158 1749 1170
rect 1583 1153 1642 1158
rect 1501 1112 1547 1124
rect 1074 1027 1290 1029
rect 1074 981 1229 1027
rect 1074 922 1105 981
rect 1219 975 1229 981
rect 1281 975 1291 1027
rect 1057 911 1105 922
rect 1584 923 1612 1153
rect 1650 1111 1719 1120
rect 1650 1077 1665 1111
rect 1699 1077 1719 1111
rect 1650 1003 1719 1077
rect 1650 969 1665 1003
rect 1699 969 1719 1003
rect 1650 952 1719 969
rect 1584 922 1630 923
rect 903 899 982 911
rect 903 863 942 899
rect 916 861 942 863
rect 936 723 942 861
rect 976 723 982 899
rect 936 711 982 723
rect 1024 899 1105 911
rect 1024 723 1030 899
rect 1064 852 1105 899
rect 1389 866 1399 918
rect 1451 914 1461 918
rect 1584 914 1661 922
rect 1451 910 1661 914
rect 1451 872 1621 910
rect 1451 866 1461 872
rect 1584 871 1621 872
rect 1064 723 1070 852
rect 1024 711 1070 723
rect 1615 734 1621 871
rect 1655 734 1661 910
rect 1615 722 1661 734
rect 1703 910 1749 922
rect 1703 734 1709 910
rect 1743 851 1749 910
rect 2066 851 2096 1205
rect 1743 758 2096 851
rect 1743 734 1749 758
rect 1703 722 1749 734
rect 1446 675 1720 681
rect 1446 674 1665 675
rect 968 664 1665 674
rect 968 630 986 664
rect 1020 641 1665 664
rect 1699 641 1720 675
rect 1020 630 1720 641
rect 968 616 1720 630
rect 541 477 741 532
rect 1263 488 1335 616
rect 1446 612 1720 616
rect 2066 489 2096 758
rect 1216 477 1335 488
rect 541 465 1335 477
rect 1615 468 1738 469
rect 1615 465 1768 468
rect 541 413 1768 465
rect 541 332 741 413
rect 839 264 885 276
rect 494 146 694 208
rect 839 146 845 264
rect 494 61 845 146
rect 494 8 694 61
rect 737 -252 765 61
rect 839 -78 845 61
rect 879 146 885 264
rect 983 272 1060 413
rect 1216 412 1768 413
rect 1216 340 1288 412
rect 1645 411 1768 412
rect 983 238 1002 272
rect 1036 238 1060 272
rect 983 230 1060 238
rect 1154 280 1201 292
rect 952 188 998 200
rect 952 146 958 188
rect 879 61 958 146
rect 879 -78 885 61
rect 952 12 958 61
rect 992 12 998 188
rect 952 0 998 12
rect 1040 188 1086 200
rect 1040 12 1046 188
rect 1080 49 1086 188
rect 1154 132 1160 280
rect 1195 264 1201 280
rect 1545 277 1591 289
rect 1545 264 1551 277
rect 1195 209 1551 264
rect 1195 132 1201 209
rect 1545 195 1551 209
rect 1585 195 1591 277
rect 1689 272 1765 411
rect 1941 289 2141 489
rect 1689 238 1709 272
rect 1743 263 1765 272
rect 1743 238 1803 263
rect 1689 237 1803 238
rect 1693 233 1803 237
rect 1697 232 1755 233
rect 1545 183 1591 195
rect 1659 188 1705 200
rect 1154 120 1201 132
rect 1659 119 1665 188
rect 1329 62 1339 119
rect 1408 118 1418 119
rect 1486 118 1589 119
rect 1634 118 1665 119
rect 1408 62 1665 118
rect 1444 61 1665 62
rect 1222 49 1232 57
rect 1080 12 1232 49
rect 1040 11 1232 12
rect 1040 0 1086 11
rect 1222 4 1232 11
rect 1285 48 1295 57
rect 1285 12 1300 48
rect 1659 12 1665 61
rect 1699 12 1705 188
rect 1285 4 1295 12
rect 1659 0 1705 12
rect 1747 188 1793 200
rect 1747 12 1753 188
rect 1787 62 1793 188
rect 2020 62 2121 289
rect 1787 27 2121 62
rect 1787 12 1793 27
rect 1747 0 1793 12
rect 1142 -28 1312 -24
rect 839 -90 885 -78
rect 987 -37 1380 -28
rect 1699 -32 1760 -31
rect 1697 -37 1760 -32
rect 987 -38 1760 -37
rect 987 -72 1002 -38
rect 1036 -72 1709 -38
rect 1743 -72 1760 -38
rect 987 -87 1760 -72
rect 987 -88 1473 -87
rect 1154 -89 1201 -88
rect 952 -252 1334 -251
rect 737 -313 1334 -252
rect 1408 -313 1419 -251
rect 737 -314 1106 -313
rect 2020 -383 2121 27
rect 1281 -384 2146 -383
rect 1220 -436 1230 -384
rect 1285 -434 2146 -384
rect 1285 -436 1951 -434
rect 2020 -436 2121 -434
<< via1 >>
rect 1397 1693 1450 1746
rect 1227 1575 1280 1628
rect 1229 975 1281 1027
rect 1399 866 1451 918
rect 1339 62 1408 119
rect 1232 4 1285 57
rect 1334 -313 1408 -251
rect 1230 -436 1285 -384
<< metal2 >>
rect 1397 1746 1450 1756
rect 1397 1683 1450 1693
rect 1227 1628 1280 1638
rect 1227 1565 1280 1575
rect 1228 1037 1280 1565
rect 1399 1564 1448 1683
rect 1228 1027 1281 1037
rect 1228 982 1229 1027
rect 1229 965 1281 975
rect 1399 918 1451 1564
rect 1399 856 1451 866
rect 1339 123 1408 129
rect 1333 119 1411 123
rect 1232 63 1285 67
rect 1231 57 1286 63
rect 1231 4 1232 57
rect 1285 4 1286 57
rect 1231 -356 1286 4
rect 1333 62 1339 119
rect 1408 62 1411 119
rect 1333 -6 1411 62
rect 1333 -37 1409 -6
rect 1333 -251 1411 -37
rect 1333 -294 1334 -251
rect 1408 -294 1411 -251
rect 1334 -323 1408 -313
rect 1230 -384 1286 -356
rect 1285 -404 1286 -384
rect 1230 -446 1285 -436
<< labels >>
flabel metal1 541 332 741 532 0 FreeSans 256 0 0 0 A
port 0 nsew
flabel metal1 404 1023 604 1223 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 1941 289 2141 489 0 FreeSans 256 0 0 0 O
port 2 nsew
flabel metal1 494 8 694 208 0 FreeSans 256 0 0 0 VSS
port 3 nsew
<< end >>
