* NGSPICE file created from inv_pex.ext - technology: sky130A

.subckt inv_pex A O VSS VDD
X0 O.t4 A.t0 VSS.t3 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 O.t0 A.t1 VDD.t5 VDD.t3 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 O.t3 A.t2 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 O.t2 A.t3 VDD.t4 VDD.t3 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 O.t5 A.t4 VDD.t2 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 O.t1 A.t5 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A.t1 A.t3 648.659
R1 A.t4 A.t5 648.644
R2 A.n0 A.t4 324.891
R3 A.n0 A.t1 324.785
R4 A.n1 A.t2 310.945
R5 A.n2 A.t0 310.073
R6 A A.n2 0.597
R7 A.n2 A.n1 0.44
R8 A.n1 A.n0 0.272
R9 VSS.n14 VSS.n9 142.811
R10 VSS.n30 VSS.n26 100.371
R11 VSS.n31 VSS.n30 81.452
R12 VSS.n15 VSS.n14 79.299
R13 VSS.n40 VSS.t1 21.252
R14 VSS.n39 VSS.t3 17.596
R15 VSS.n32 VSS.n31 15
R16 VSS.n33 VSS.n32 15
R17 VSS.n25 VSS.n15 14.711
R18 VSS.n23 VSS.n22 14.102
R19 VSS.n38 VSS.n37 13.653
R20 VSS.n38 VSS.n36 2.44
R21 VSS.n26 VSS.n25 0.967
R22 VSS VSS.n40 0.208
R23 VSS.n40 VSS.n39 0.163
R24 VSS.n25 VSS.n24 0.146
R25 VSS.n24 VSS.n23 0.138
R26 VSS.n6 VSS.n5 0.062
R27 VSS.n7 VSS.n6 0.062
R28 VSS.n26 VSS.n7 0.054
R29 VSS.n39 VSS.n38 0.026
R30 VSS.n23 VSS.n21 0.009
R31 VSS.n3 VSS.n2 0.003
R32 VSS.n4 VSS.n3 0.003
R33 VSS.n14 VSS.n13 0.003
R34 VSS.n13 VSS.t0 0.003
R35 VSS.n11 VSS.n10 0.003
R36 VSS.n30 VSS.n29 0.003
R37 VSS.n29 VSS.t2 0.003
R38 VSS.t2 VSS.n28 0.003
R39 VSS.n28 VSS.n27 0.003
R40 VSS.n20 VSS.n17 0.002
R41 VSS.n20 VSS.n19 0.002
R42 VSS.n5 VSS.n1 0.002
R43 VSS.n12 VSS.n11 0.002
R44 VSS.n34 VSS.n33 0.002
R45 VSS.n17 VSS.n16 0.002
R46 VSS.n19 VSS.n18 0.002
R47 VSS.n1 VSS.n0 0.002
R48 VSS.n36 VSS.n35 0.002
R49 VSS.n35 VSS.n34 0.002
R50 VSS.t0 VSS.n12 0.001
R51 VSS.n9 VSS.n8 0.001
R52 VSS.n5 VSS.n4 0.001
R53 VSS.n21 VSS.n20 0.001
R54 O.n1 O.t2 29.729
R55 O.n2 O.t1 29.072
R56 O.n3 O.t5 29.072
R57 O.n1 O.t0 29.062
R58 O.n0 O.t4 21.547
R59 O.n0 O.t3 18.392
R60 O.n2 O.n1 7.248
R61 O.n3 O.n2 1.475
R62 O O.n3 1.245
R63 O O.n0 0.303
R64 VDD.n15 VDD.n14 99.394
R65 VDD.n6 VDD.n5 94.207
R66 VDD.n20 VDD.n17 83.233
R67 VDD.n22 VDD.t1 31.277
R68 VDD.n0 VDD.t5 29.922
R69 VDD.n0 VDD.t4 29.596
R70 VDD.n22 VDD.t2 28.803
R71 VDD.n12 VDD.n10 22.354
R72 VDD.n10 VDD.n8 7.569
R73 VDD.n23 VDD.n22 7.452
R74 VDD.n10 VDD.n9 4.546
R75 VDD.n8 VDD.n7 1.322
R76 VDD.n12 VDD.n11 1.288
R77 VDD VDD.n23 0.285
R78 VDD.n23 VDD.n21 0.199
R79 VDD.n21 VDD.n0 0.148
R80 VDD.n7 VDD.n6 0.084
R81 VDD.n21 VDD.n20 0.069
R82 VDD.n6 VDD.n2 0.009
R83 VDD.n2 VDD.n1 0.008
R84 VDD.n14 VDD.n13 0.008
R85 VDD.n13 VDD.n12 0.008
R86 VDD.n17 VDD.t3 0.004
R87 VDD.n20 VDD.n19 0.003
R88 VDD.n19 VDD.n18 0.003
R89 VDD.n4 VDD.n3 0.003
R90 VDD.n5 VDD.t0 0.003
R91 VDD.t0 VDD.n4 0.003
R92 VDD.n16 VDD.n15 0.003
R93 VDD.t3 VDD.n16 0.003
C0 VDD A 3.02fF
C1 O VDD 3.71fF
C2 O A 1.63fF
.ends

