magic
tech sky130A
magscale 1 2
timestamp 1659038648
<< pwell >>
rect -307 -1378 307 1378
<< psubdiff >>
rect -271 1308 -175 1342
rect 175 1308 271 1342
rect -271 1246 -237 1308
rect 237 1246 271 1308
rect -271 -1308 -237 -1246
rect 237 -1308 271 -1246
rect -271 -1342 -175 -1308
rect 175 -1342 271 -1308
<< psubdiffcont >>
rect -175 1308 175 1342
rect -271 -1246 -237 1246
rect 237 -1246 271 1246
rect -175 -1342 175 -1308
<< xpolycontact >>
rect -141 780 141 1212
rect -141 -1212 141 -780
<< xpolyres >>
rect -141 -780 141 780
<< locali >>
rect -271 1308 -175 1342
rect 175 1308 271 1342
rect -271 1246 -237 1308
rect 237 1246 271 1308
rect -271 -1308 -237 -1246
rect 237 -1308 271 -1246
rect -271 -1342 -175 -1308
rect 175 -1342 271 -1308
<< viali >>
rect -125 797 125 1194
rect -125 -1194 125 -797
<< metal1 >>
rect -131 1194 131 1206
rect -131 797 -125 1194
rect 125 797 131 1194
rect -131 785 131 797
rect -131 -797 131 -785
rect -131 -1194 -125 -797
rect 125 -1194 131 -797
rect -131 -1206 131 -1194
<< res1p41 >>
rect -143 -782 143 782
<< properties >>
string FIXED_BBOX -254 -1325 254 1325
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 7.8 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 11.091k dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
