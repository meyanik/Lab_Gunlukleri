magic
tech sky130A
magscale 1 2
timestamp 1658993734
<< nwell >>
rect -496 -2573 496 2573
<< pmoslvt >>
rect -300 1354 300 2354
rect -300 118 300 1118
rect -300 -1118 300 -118
rect -300 -2354 300 -1354
<< pdiff >>
rect -358 2342 -300 2354
rect -358 1366 -346 2342
rect -312 1366 -300 2342
rect -358 1354 -300 1366
rect 300 2342 358 2354
rect 300 1366 312 2342
rect 346 1366 358 2342
rect 300 1354 358 1366
rect -358 1106 -300 1118
rect -358 130 -346 1106
rect -312 130 -300 1106
rect -358 118 -300 130
rect 300 1106 358 1118
rect 300 130 312 1106
rect 346 130 358 1106
rect 300 118 358 130
rect -358 -130 -300 -118
rect -358 -1106 -346 -130
rect -312 -1106 -300 -130
rect -358 -1118 -300 -1106
rect 300 -130 358 -118
rect 300 -1106 312 -130
rect 346 -1106 358 -130
rect 300 -1118 358 -1106
rect -358 -1366 -300 -1354
rect -358 -2342 -346 -1366
rect -312 -2342 -300 -1366
rect -358 -2354 -300 -2342
rect 300 -1366 358 -1354
rect 300 -2342 312 -1366
rect 346 -2342 358 -1366
rect 300 -2354 358 -2342
<< pdiffc >>
rect -346 1366 -312 2342
rect 312 1366 346 2342
rect -346 130 -312 1106
rect 312 130 346 1106
rect -346 -1106 -312 -130
rect 312 -1106 346 -130
rect -346 -2342 -312 -1366
rect 312 -2342 346 -1366
<< nsubdiff >>
rect -460 2503 -364 2537
rect 364 2503 460 2537
rect -460 2441 -426 2503
rect 426 2441 460 2503
rect -460 -2503 -426 -2441
rect 426 -2503 460 -2441
rect -460 -2537 -364 -2503
rect 364 -2537 460 -2503
<< nsubdiffcont >>
rect -364 2503 364 2537
rect -460 -2441 -426 2441
rect 426 -2441 460 2441
rect -364 -2537 364 -2503
<< poly >>
rect -300 2435 300 2451
rect -300 2401 -284 2435
rect 284 2401 300 2435
rect -300 2354 300 2401
rect -300 1307 300 1354
rect -300 1273 -284 1307
rect 284 1273 300 1307
rect -300 1257 300 1273
rect -300 1199 300 1215
rect -300 1165 -284 1199
rect 284 1165 300 1199
rect -300 1118 300 1165
rect -300 71 300 118
rect -300 37 -284 71
rect 284 37 300 71
rect -300 21 300 37
rect -300 -37 300 -21
rect -300 -71 -284 -37
rect 284 -71 300 -37
rect -300 -118 300 -71
rect -300 -1165 300 -1118
rect -300 -1199 -284 -1165
rect 284 -1199 300 -1165
rect -300 -1215 300 -1199
rect -300 -1273 300 -1257
rect -300 -1307 -284 -1273
rect 284 -1307 300 -1273
rect -300 -1354 300 -1307
rect -300 -2401 300 -2354
rect -300 -2435 -284 -2401
rect 284 -2435 300 -2401
rect -300 -2451 300 -2435
<< polycont >>
rect -284 2401 284 2435
rect -284 1273 284 1307
rect -284 1165 284 1199
rect -284 37 284 71
rect -284 -71 284 -37
rect -284 -1199 284 -1165
rect -284 -1307 284 -1273
rect -284 -2435 284 -2401
<< locali >>
rect -460 2503 -364 2537
rect 364 2503 460 2537
rect -460 2441 -426 2503
rect 426 2441 460 2503
rect -300 2401 -284 2435
rect 284 2401 300 2435
rect -346 2342 -312 2358
rect -346 1350 -312 1366
rect 312 2342 346 2358
rect 312 1350 346 1366
rect -300 1273 -284 1307
rect 284 1273 300 1307
rect -300 1165 -284 1199
rect 284 1165 300 1199
rect -346 1106 -312 1122
rect -346 114 -312 130
rect 312 1106 346 1122
rect 312 114 346 130
rect -300 37 -284 71
rect 284 37 300 71
rect -300 -71 -284 -37
rect 284 -71 300 -37
rect -346 -130 -312 -114
rect -346 -1122 -312 -1106
rect 312 -130 346 -114
rect 312 -1122 346 -1106
rect -300 -1199 -284 -1165
rect 284 -1199 300 -1165
rect -300 -1307 -284 -1273
rect 284 -1307 300 -1273
rect -346 -1366 -312 -1350
rect -346 -2358 -312 -2342
rect 312 -1366 346 -1350
rect 312 -2358 346 -2342
rect -300 -2435 -284 -2401
rect 284 -2435 300 -2401
rect -460 -2503 -426 -2441
rect 426 -2503 460 -2441
rect -460 -2537 -364 -2503
rect 364 -2537 460 -2503
<< viali >>
rect -284 2401 284 2435
rect -346 1366 -312 2342
rect 312 1366 346 2342
rect -284 1273 284 1307
rect -284 1165 284 1199
rect -346 130 -312 1106
rect 312 130 346 1106
rect -284 37 284 71
rect -284 -71 284 -37
rect -346 -1106 -312 -130
rect 312 -1106 346 -130
rect -284 -1199 284 -1165
rect -284 -1307 284 -1273
rect -346 -2342 -312 -1366
rect 312 -2342 346 -1366
rect -284 -2435 284 -2401
<< metal1 >>
rect -296 2435 296 2441
rect -296 2401 -284 2435
rect 284 2401 296 2435
rect -296 2395 296 2401
rect -352 2342 -306 2354
rect -352 1366 -346 2342
rect -312 1366 -306 2342
rect -352 1354 -306 1366
rect 306 2342 352 2354
rect 306 1366 312 2342
rect 346 1366 352 2342
rect 306 1354 352 1366
rect -296 1307 296 1313
rect -296 1273 -284 1307
rect 284 1273 296 1307
rect -296 1267 296 1273
rect -296 1199 296 1205
rect -296 1165 -284 1199
rect 284 1165 296 1199
rect -296 1159 296 1165
rect -352 1106 -306 1118
rect -352 130 -346 1106
rect -312 130 -306 1106
rect -352 118 -306 130
rect 306 1106 352 1118
rect 306 130 312 1106
rect 346 130 352 1106
rect 306 118 352 130
rect -296 71 296 77
rect -296 37 -284 71
rect 284 37 296 71
rect -296 31 296 37
rect -296 -37 296 -31
rect -296 -71 -284 -37
rect 284 -71 296 -37
rect -296 -77 296 -71
rect -352 -130 -306 -118
rect -352 -1106 -346 -130
rect -312 -1106 -306 -130
rect -352 -1118 -306 -1106
rect 306 -130 352 -118
rect 306 -1106 312 -130
rect 346 -1106 352 -130
rect 306 -1118 352 -1106
rect -296 -1165 296 -1159
rect -296 -1199 -284 -1165
rect 284 -1199 296 -1165
rect -296 -1205 296 -1199
rect -296 -1273 296 -1267
rect -296 -1307 -284 -1273
rect 284 -1307 296 -1273
rect -296 -1313 296 -1307
rect -352 -1366 -306 -1354
rect -352 -2342 -346 -1366
rect -312 -2342 -306 -1366
rect -352 -2354 -306 -2342
rect 306 -1366 352 -1354
rect 306 -2342 312 -1366
rect 346 -2342 352 -1366
rect 306 -2354 352 -2342
rect -296 -2401 296 -2395
rect -296 -2435 -284 -2401
rect 284 -2435 296 -2401
rect -296 -2441 296 -2435
<< properties >>
string FIXED_BBOX -443 -2520 443 2520
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 5.0 l 3.0 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
