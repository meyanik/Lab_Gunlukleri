magic
tech sky130A
magscale 1 2
timestamp 1659200772
<< nwell >>
rect -12938 8167 -12905 8247
rect -12938 8163 -12880 8167
rect -15661 8099 -15624 8105
rect -15661 7957 -15630 7961
rect -15661 7951 -15624 7957
rect -12938 7884 -12910 8163
rect -12369 7901 -12349 8163
rect -11492 7909 -11464 8158
rect -12913 7804 -12910 7884
<< pwell >>
rect -19328 5944 -18927 5947
rect -20918 5893 -20844 5901
rect -19584 4669 -19556 4900
rect -19447 4803 -19439 4807
rect -19447 4716 -19419 4803
rect -16981 4730 -16953 4799
rect -14289 4794 -14107 5104
rect -19584 4640 -19548 4669
rect -17285 4112 -17106 4140
rect -18708 3539 -18680 3540
rect -18837 3512 -18680 3539
rect -16841 3523 -16812 3680
rect -16164 3525 -16135 3682
rect -15490 3530 -15461 3687
rect -14791 3526 -14762 3683
rect -18877 3511 -18680 3512
<< viali >>
rect -18042 7711 -18007 8083
rect -17663 7710 -17628 8082
rect -16776 7706 -16742 8067
rect -16416 7706 -16382 8067
rect -15530 7706 -15496 8067
rect -15170 7706 -15136 8067
rect -14284 7707 -14250 8069
rect -13922 7708 -13888 8070
rect -12836 7708 -12802 8070
rect -12476 7710 -12442 8072
rect -13696 5960 -13196 5994
rect -13696 5868 -13196 5902
rect -13696 5360 -13196 5394
rect -13696 5254 -13196 5288
rect -14492 4590 -13951 4691
rect -13694 4590 -13153 4691
rect -12896 4590 -12355 4691
rect -12099 4590 -11456 4691
rect -14431 4456 -14037 4528
rect -13609 4456 -13239 4528
rect -12811 4456 -12441 4528
rect -12013 4527 -11643 4528
rect -12013 4456 -11619 4527
rect -14431 4110 -14359 4456
rect -11691 4110 -11619 4456
rect -11557 3947 -11456 4590
rect -20155 3717 -20083 3781
rect -20331 3645 -20083 3717
rect -20021 3482 -19920 3781
rect -14439 3384 -14367 3730
rect -11699 3384 -11627 3729
rect -14439 3312 -14045 3384
rect -13617 3312 -13247 3384
rect -12819 3312 -12449 3384
rect -12021 3312 -11627 3384
rect -11565 3250 -11464 3893
rect -14501 3149 -13959 3250
rect -13703 3149 -13161 3250
rect -12905 3149 -12363 3250
rect -12107 3149 -11464 3250
rect -20511 960 -20477 1053
rect -20423 960 -20389 1053
<< metal1 >>
rect -20274 9467 -20264 9519
rect -20212 9505 -20202 9519
rect -19086 9505 -19076 9517
rect -20212 9477 -19076 9505
rect -20212 9467 -20202 9477
rect -19086 9465 -19076 9477
rect -19024 9508 -19014 9517
rect -17802 9508 -17792 9511
rect -19024 9480 -17792 9508
rect -19024 9465 -19014 9480
rect -17802 9459 -17792 9480
rect -17740 9502 -17730 9511
rect -16539 9502 -16529 9512
rect -17740 9474 -16529 9502
rect -17740 9459 -17730 9474
rect -16539 9460 -16529 9474
rect -16477 9502 -16467 9512
rect -15278 9502 -15268 9514
rect -16477 9474 -15268 9502
rect -16477 9460 -16467 9474
rect -15278 9462 -15268 9474
rect -15216 9502 -15206 9514
rect -14027 9502 -14017 9512
rect -15216 9474 -14017 9502
rect -15216 9462 -15206 9474
rect -14027 9460 -14017 9474
rect -13965 9502 -13955 9512
rect -12576 9502 -12566 9511
rect -13965 9474 -12566 9502
rect -13965 9460 -13955 9474
rect -12576 9459 -12566 9474
rect -12514 9459 -12504 9511
rect -17950 9392 -17942 9444
rect -17890 9430 -17880 9444
rect -17890 9425 -17879 9430
rect -16688 9425 -16678 9440
rect -17890 9396 -16678 9425
rect -17890 9392 -17880 9396
rect -16688 9388 -16678 9396
rect -16626 9388 -16616 9440
rect -12772 9370 -12762 9422
rect -12710 9416 -12700 9422
rect -11324 9416 -11314 9429
rect -12710 9388 -11314 9416
rect -12710 9370 -12700 9388
rect -11324 9377 -11314 9388
rect -11262 9377 -11252 9429
rect -12772 9115 -12762 9128
rect -12928 9086 -12762 9115
rect -16688 9065 -16678 9076
rect -16864 9031 -16678 9065
rect -16688 9024 -16678 9031
rect -16626 9024 -16616 9076
rect -12772 9074 -12762 9086
rect -12709 9074 -12699 9128
rect -20273 8920 -20263 8972
rect -20211 8965 -20201 8972
rect -19086 8966 -19076 9018
rect -19024 9010 -19014 9018
rect -19024 8975 -18798 9010
rect -17953 8981 -17943 8988
rect -19024 8966 -19014 8975
rect -20211 8930 -20035 8965
rect -18124 8940 -17943 8981
rect -17953 8936 -17943 8940
rect -17891 8936 -17881 8988
rect -20211 8920 -20201 8930
rect -16541 8915 -16531 8967
rect -16479 8959 -16469 8967
rect -16479 8924 -16274 8959
rect -16479 8915 -16469 8924
rect -15278 8909 -15268 8961
rect -15216 8954 -15206 8961
rect -15216 8918 -15043 8954
rect -15216 8909 -15206 8918
rect -14026 8909 -14016 8961
rect -13964 8953 -13954 8961
rect -13964 8917 -13807 8953
rect -13964 8909 -13954 8917
rect -12577 8908 -12567 8960
rect -12515 8953 -12505 8960
rect -12515 8917 -12360 8953
rect -12515 8908 -12505 8917
rect -11324 8786 -11314 8794
rect -11478 8751 -11314 8786
rect -11324 8742 -11314 8751
rect -11262 8742 -11252 8794
rect -17802 8550 -17792 8602
rect -17740 8595 -17730 8602
rect -17740 8554 -17542 8595
rect -17740 8550 -17730 8554
rect -19205 8230 -19195 8238
rect -19377 8196 -19195 8230
rect -19205 8186 -19195 8196
rect -19143 8186 -19133 8238
rect -20922 7875 -20884 8161
rect -20774 7985 -20742 8084
rect -20634 7888 -20596 8174
rect -18823 8096 -18795 8192
rect -19575 8073 -19553 8075
rect -20350 7751 -20340 7803
rect -20288 7792 -20278 7803
rect -19777 7792 -19767 7805
rect -20288 7763 -19767 7792
rect -20288 7751 -20278 7763
rect -19777 7753 -19767 7763
rect -19715 7753 -19705 7805
rect -19575 7520 -19546 8073
rect -19438 8067 -18752 8096
rect -18823 7873 -18795 8067
rect -18432 7975 -18394 8074
rect -18142 7882 -18108 8182
rect -18048 8083 -18001 8095
rect -18048 7711 -18042 8083
rect -18007 7875 -18001 8083
rect -17669 8082 -17622 8094
rect -17669 7875 -17663 8082
rect -18007 7846 -17663 7875
rect -18007 7711 -18001 7846
rect -18048 7699 -18001 7711
rect -17669 7710 -17663 7846
rect -17628 7710 -17622 8082
rect -17561 7880 -17531 8204
rect -17177 7982 -17140 8077
rect -16877 7868 -16847 8192
rect -15633 8105 -15604 8158
rect -14387 8105 -14358 8158
rect -15661 8100 -15604 8105
rect -15665 8099 -15604 8100
rect -16782 8067 -16736 8079
rect -17669 7698 -17622 7710
rect -16782 7706 -16776 8067
rect -16742 7904 -16736 8067
rect -16422 8067 -16376 8079
rect -16422 7904 -16416 8067
rect -16742 7875 -16416 7904
rect -16742 7706 -16736 7875
rect -16782 7694 -16736 7706
rect -16422 7706 -16416 7875
rect -16382 7706 -16376 8067
rect -15667 8059 -15604 8099
rect -15632 7997 -15604 8059
rect -15667 7961 -15604 7997
rect -15665 7960 -15604 7961
rect -15661 7951 -15604 7960
rect -15633 7894 -15604 7951
rect -15536 8067 -15490 8079
rect -16422 7694 -16376 7706
rect -15536 7706 -15530 8067
rect -15496 7915 -15490 8067
rect -15176 8067 -15130 8079
rect -15176 7915 -15170 8067
rect -15496 7886 -15170 7915
rect -15496 7706 -15490 7886
rect -15536 7694 -15490 7706
rect -15176 7706 -15170 7886
rect -15136 7706 -15130 8067
rect -14427 8057 -14358 8105
rect -14387 7997 -14358 8057
rect -14436 7951 -14358 7997
rect -14387 7888 -14358 7951
rect -14290 8069 -14244 8081
rect -15176 7694 -15130 7706
rect -14290 7707 -14284 8069
rect -14250 7895 -14244 8069
rect -13928 8070 -13882 8082
rect -13928 7895 -13922 8070
rect -14250 7866 -13922 7895
rect -14250 7707 -14244 7866
rect -14290 7695 -14244 7707
rect -13928 7708 -13922 7866
rect -13888 7708 -13882 8070
rect -13819 7857 -13786 8220
rect -12938 8163 -12905 8247
rect -13454 8060 -13446 8074
rect -13455 7996 -13426 8060
rect -13454 7979 -13446 7996
rect -12938 7884 -12910 8163
rect -12369 8150 -12349 8163
rect -11492 8153 -11464 8158
rect -12933 7800 -12910 7884
rect -12842 8070 -12796 8082
rect -13928 7696 -13882 7708
rect -12842 7708 -12836 8070
rect -12802 7930 -12796 8070
rect -12482 8072 -12436 8084
rect -12482 7930 -12476 8072
rect -12802 7901 -12476 7930
rect -12802 7708 -12796 7901
rect -12842 7696 -12796 7708
rect -12482 7710 -12476 7901
rect -12442 7710 -12436 8072
rect -12369 7901 -12341 8150
rect -11876 7993 -11846 8062
rect -11492 7909 -11463 8153
rect -11491 7904 -11463 7909
rect -12482 7698 -12436 7710
rect -20349 7367 -20339 7419
rect -20287 7404 -20277 7419
rect -20287 7375 -20042 7404
rect -20287 7367 -20277 7375
rect -21165 6927 -21155 6981
rect -21102 6967 -21092 6981
rect -20456 6976 -20446 6989
rect -21102 6938 -20899 6967
rect -20625 6946 -20446 6976
rect -21102 6927 -21092 6938
rect -20456 6935 -20446 6946
rect -20393 6935 -20383 6989
rect -20371 6862 -20361 6875
rect -20674 6832 -20361 6862
rect -20371 6821 -20361 6832
rect -20308 6821 -20298 6875
rect -15313 6861 -15303 6872
rect -18220 6850 -17466 6859
rect -18220 6828 -17449 6850
rect -16930 6831 -16197 6861
rect -15692 6831 -15303 6861
rect -15313 6820 -15303 6831
rect -15251 6861 -15241 6872
rect -15251 6831 -14959 6861
rect -14435 6831 -13742 6861
rect -12987 6831 -12294 6861
rect -15251 6820 -15241 6831
rect -19215 6583 -19205 6594
rect -19370 6553 -19205 6583
rect -19215 6540 -19205 6553
rect -19152 6540 -19142 6594
rect -21167 6368 -21157 6423
rect -21102 6404 -21092 6423
rect -21102 6375 -20000 6404
rect -21102 6368 -21092 6375
rect -20370 6161 -20362 6216
rect -20309 6199 -20299 6216
rect -19216 6199 -19206 6214
rect -20309 6170 -19206 6199
rect -20309 6161 -20299 6170
rect -19216 6160 -19206 6170
rect -19153 6160 -19143 6214
rect -16689 6133 -16679 6147
rect -20441 6132 -20267 6133
rect -17865 6132 -16679 6133
rect -20441 6130 -16679 6132
rect -20457 6074 -20447 6130
rect -20393 6103 -16679 6130
rect -20393 6074 -20383 6103
rect -18566 5947 -18518 6103
rect -16689 6093 -16679 6103
rect -16626 6093 -16616 6147
rect -14793 6137 -14238 6339
rect -19328 5944 -18927 5947
rect -20918 5894 -20844 5901
rect -20651 5900 -20445 5901
rect -20371 5900 -20361 5919
rect -20918 5873 -20838 5894
rect -20651 5873 -20361 5900
rect -20918 5834 -20882 5873
rect -20516 5872 -20361 5873
rect -20371 5864 -20361 5872
rect -20308 5864 -20298 5919
rect -19575 5904 -19517 5944
rect -19335 5919 -18926 5944
rect -18738 5919 -17544 5947
rect -19575 5844 -19547 5904
rect -18984 5859 -18956 5919
rect -18566 5918 -18518 5919
rect -18392 5869 -18364 5919
rect -17800 5869 -17772 5919
rect -16872 5916 -16383 5944
rect -16196 5916 -15011 5944
rect -14792 5775 -14764 6137
rect -13708 5994 -13184 6000
rect -13708 5960 -13696 5994
rect -13196 5960 -13184 5994
rect -13708 5954 -13184 5960
rect -13545 5908 -13421 5954
rect -13708 5902 -13184 5908
rect -13708 5868 -13696 5902
rect -13196 5868 -13184 5902
rect -13708 5862 -13184 5868
rect -12308 5737 -12127 6178
rect -20581 5112 -20266 5146
rect -14293 5106 -14112 5547
rect -13708 5394 -13184 5400
rect -13708 5360 -13696 5394
rect -13196 5360 -13184 5394
rect -13708 5354 -13184 5360
rect -13541 5294 -13417 5354
rect -13708 5288 -13184 5294
rect -13708 5254 -13696 5288
rect -13196 5254 -13184 5288
rect -13708 5248 -13184 5254
rect -12290 5106 -12109 5547
rect -19584 4900 -19566 4905
rect -19584 4669 -19556 4900
rect -19447 4803 -19439 4807
rect -19447 4716 -19419 4803
rect -19584 4640 -19548 4669
rect -19300 4652 -19272 4888
rect -18985 4645 -18957 4881
rect -18846 4731 -18818 4795
rect -18708 4646 -18680 4882
rect -18392 4643 -18364 4878
rect -18258 4718 -18230 4819
rect -18116 4646 -18088 4881
rect -17800 4644 -17772 4879
rect -17666 4712 -17638 4813
rect -17524 4642 -17496 4877
rect -17118 4642 -17090 4876
rect -16981 4730 -16953 4799
rect -16842 4649 -16814 4893
rect -16444 4641 -16416 4882
rect -16309 4728 -16281 4797
rect -16168 4636 -16140 4880
rect -15766 4641 -15738 4880
rect -15633 4730 -15605 4799
rect -15490 4640 -15462 4879
rect -15068 4643 -15040 4882
rect -14932 4731 -14904 4800
rect -14792 4642 -14764 4881
rect -14289 4834 -14107 5104
rect -14289 4794 -13837 4834
rect -14504 4691 -13939 4697
rect -14504 4590 -14492 4691
rect -13951 4590 -13939 4691
rect -14504 4584 -13939 4590
rect -19799 4548 -19789 4561
rect -19938 4520 -19789 4548
rect -19799 4506 -19789 4520
rect -19736 4506 -19726 4561
rect -14437 4534 -14353 4540
rect -14265 4534 -14226 4584
rect -14437 4528 -14025 4534
rect -20280 4425 -20248 4487
rect -20280 4397 -20167 4425
rect -17349 4098 -17339 4153
rect -17286 4140 -17276 4153
rect -17286 4138 -17106 4140
rect -17286 4112 -17101 4138
rect -16678 4129 -16668 4185
rect -16614 4174 -16604 4185
rect -16614 4146 -16431 4174
rect -16614 4129 -16604 4146
rect -15997 4136 -15987 4191
rect -15933 4182 -15923 4191
rect -15933 4154 -15747 4182
rect -15933 4136 -15923 4154
rect -15314 4138 -15304 4194
rect -15250 4187 -15240 4194
rect -15250 4159 -15064 4187
rect -15250 4138 -15240 4159
rect -17286 4098 -17276 4112
rect -14437 4110 -14431 4528
rect -14037 4456 -14025 4528
rect -14359 4450 -14025 4456
rect -14359 4110 -14353 4450
rect -13911 4333 -13838 4794
rect -11563 4697 -11450 4703
rect -13706 4691 -13141 4697
rect -13706 4590 -13694 4691
rect -13153 4661 -13141 4691
rect -12908 4691 -12343 4697
rect -12908 4661 -12896 4691
rect -13153 4615 -12896 4661
rect -13153 4590 -13141 4615
rect -13706 4584 -13141 4590
rect -12908 4590 -12896 4615
rect -12355 4663 -12343 4691
rect -12111 4691 -11450 4697
rect -12111 4663 -12099 4691
rect -12355 4617 -12099 4663
rect -12355 4590 -12343 4617
rect -12908 4584 -12343 4590
rect -12111 4590 -12099 4617
rect -12111 4584 -11557 4590
rect -13448 4534 -13409 4584
rect -12642 4534 -12603 4584
rect -11846 4534 -11807 4584
rect -11697 4534 -11613 4539
rect -13621 4528 -13227 4534
rect -13621 4456 -13609 4528
rect -13239 4456 -13227 4528
rect -13621 4450 -13227 4456
rect -12823 4528 -12429 4534
rect -12823 4456 -12811 4528
rect -12441 4456 -12429 4528
rect -12823 4450 -12429 4456
rect -12025 4528 -11613 4534
rect -12025 4456 -12013 4528
rect -11643 4527 -11613 4528
rect -12025 4450 -11691 4456
rect -14158 4293 -13450 4333
rect -13364 4300 -12656 4340
rect -12571 4301 -11863 4341
rect -13911 4291 -13838 4293
rect -14437 4098 -14353 4110
rect -19881 3877 -19871 3886
rect -20227 3840 -19871 3877
rect -19881 3831 -19871 3840
rect -19818 3831 -19808 3886
rect -20161 3781 -19914 3793
rect -20161 3723 -20155 3781
rect -20343 3717 -20155 3723
rect -20343 3645 -20331 3717
rect -20083 3645 -20021 3781
rect -20343 3639 -20021 3645
rect -20084 3638 -20021 3639
rect -20027 3482 -20021 3638
rect -19920 3482 -19914 3781
rect -14421 3742 -14371 4098
rect -14445 3730 -14361 3742
rect -19883 3502 -19873 3557
rect -19820 3539 -19810 3557
rect -19300 3539 -19272 3669
rect -18708 3539 -18680 3677
rect -17526 3654 -17496 3662
rect -17524 3539 -17496 3654
rect -19820 3511 -17496 3539
rect -16841 3538 -16812 3680
rect -16164 3538 -16135 3682
rect -15490 3538 -15461 3687
rect -14791 3538 -14762 3683
rect -19820 3502 -19810 3511
rect -16845 3510 -14735 3538
rect -20027 3470 -19914 3482
rect -17349 3403 -17339 3459
rect -17286 3434 -17276 3459
rect -16676 3434 -16666 3456
rect -17286 3403 -16666 3434
rect -16676 3400 -16666 3403
rect -16612 3434 -16602 3456
rect -15994 3434 -15984 3459
rect -16612 3404 -15984 3434
rect -15931 3434 -15921 3459
rect -15314 3434 -15304 3458
rect -15931 3404 -15304 3434
rect -16612 3403 -15304 3404
rect -15251 3403 -15241 3458
rect -16612 3400 -16602 3403
rect -14445 3312 -14439 3730
rect -14367 3390 -14361 3730
rect -14246 3595 -14206 4257
rect -11697 4110 -11691 4450
rect -11619 4110 -11613 4527
rect -11697 4098 -11613 4110
rect -11563 3947 -11557 4584
rect -11456 3947 -11450 4691
rect -11563 3935 -11450 3947
rect -11549 3905 -11465 3935
rect -11571 3893 -11458 3905
rect -11705 3729 -11621 3741
rect -14175 3503 -13467 3543
rect -13380 3501 -12672 3541
rect -12586 3507 -11878 3547
rect -11705 3390 -11699 3729
rect -14367 3384 -14033 3390
rect -14045 3312 -14033 3384
rect -14445 3306 -14033 3312
rect -13629 3384 -13235 3390
rect -13629 3312 -13617 3384
rect -13247 3312 -13235 3384
rect -13629 3306 -13235 3312
rect -12831 3384 -12437 3390
rect -12831 3312 -12819 3384
rect -12449 3312 -12437 3384
rect -12831 3306 -12437 3312
rect -12033 3384 -11699 3390
rect -12033 3312 -12021 3384
rect -11627 3312 -11621 3729
rect -12033 3306 -11621 3312
rect -14445 3300 -14361 3306
rect -14247 3256 -14208 3306
rect -13454 3256 -13415 3306
rect -12658 3256 -12619 3306
rect -11856 3256 -11817 3306
rect -11705 3300 -11621 3306
rect -11571 3256 -11565 3893
rect -14513 3250 -13947 3256
rect -14513 3149 -14501 3250
rect -13959 3222 -13947 3250
rect -13715 3250 -13149 3256
rect -13715 3222 -13703 3250
rect -13959 3176 -13703 3222
rect -13959 3149 -13947 3176
rect -14513 3143 -13947 3149
rect -13715 3149 -13703 3176
rect -13161 3222 -13149 3250
rect -12917 3250 -12351 3256
rect -12917 3222 -12905 3250
rect -13161 3176 -12905 3222
rect -13161 3149 -13149 3176
rect -13715 3143 -13149 3149
rect -12917 3149 -12905 3176
rect -12363 3222 -12351 3250
rect -12119 3250 -11565 3256
rect -11464 3256 -11458 3893
rect -12119 3222 -12107 3250
rect -12363 3176 -12107 3222
rect -12363 3149 -12351 3176
rect -12917 3143 -12351 3149
rect -12119 3149 -12107 3176
rect -11464 3149 -11452 3256
rect -12119 3143 -11452 3149
rect -11571 3137 -11458 3143
rect -20517 1053 -20471 1065
rect -20517 960 -20511 1053
rect -20477 960 -20471 1053
rect -20517 948 -20471 960
rect -20429 1053 -20383 1065
rect -20429 960 -20423 1053
rect -20389 960 -20383 1053
rect -20429 948 -20383 960
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
<< via1 >>
rect -20264 9467 -20212 9519
rect -19076 9465 -19024 9517
rect -17792 9459 -17740 9511
rect -16529 9460 -16477 9512
rect -15268 9462 -15216 9514
rect -14017 9460 -13965 9512
rect -12566 9459 -12514 9511
rect -17942 9392 -17890 9444
rect -16678 9388 -16626 9440
rect -12762 9370 -12710 9422
rect -11314 9377 -11262 9429
rect -16678 9024 -16626 9076
rect -12762 9074 -12709 9128
rect -20263 8920 -20211 8972
rect -19076 8966 -19024 9018
rect -17943 8936 -17891 8988
rect -16531 8915 -16479 8967
rect -15268 8909 -15216 8961
rect -14016 8909 -13964 8961
rect -12567 8908 -12515 8960
rect -11314 8742 -11262 8794
rect -17792 8550 -17740 8602
rect -19195 8186 -19143 8238
rect -20340 7751 -20288 7803
rect -19767 7753 -19715 7805
rect -20339 7367 -20287 7419
rect -21155 6927 -21102 6981
rect -20446 6935 -20393 6989
rect -20361 6821 -20308 6875
rect -15303 6820 -15251 6872
rect -19205 6540 -19152 6594
rect -21157 6368 -21102 6423
rect -20362 6161 -20309 6216
rect -19206 6160 -19153 6214
rect -20447 6074 -20393 6130
rect -16679 6093 -16626 6147
rect -20361 5864 -20308 5919
rect -19789 4506 -19736 4561
rect -17339 4098 -17286 4153
rect -16668 4129 -16614 4185
rect -15987 4136 -15933 4191
rect -15304 4138 -15250 4194
rect -19871 3831 -19818 3886
rect -19873 3502 -19820 3557
rect -17339 3403 -17286 3459
rect -16666 3400 -16612 3456
rect -15984 3404 -15931 3459
rect -15304 3403 -15251 3458
<< metal2 >>
rect -20264 9519 -20212 9529
rect -20264 9457 -20212 9467
rect -19076 9517 -19024 9527
rect -17792 9511 -17740 9521
rect -20259 9406 -20213 9457
rect -19076 9455 -19024 9465
rect -20259 8982 -20214 9406
rect -19073 9028 -19027 9455
rect -17943 9444 -17889 9511
rect -17943 9392 -17942 9444
rect -17890 9392 -17889 9444
rect -19076 9018 -19024 9028
rect -20263 8972 -20211 8982
rect -19076 8956 -19024 8966
rect -17943 8988 -17889 9392
rect -17891 8936 -17889 8988
rect -17943 8925 -17889 8936
rect -17793 9459 -17792 9487
rect -16529 9512 -16477 9522
rect -17740 9459 -17739 9487
rect -20263 8910 -20211 8920
rect -17793 8602 -17739 9459
rect -16529 9450 -16477 9460
rect -15268 9514 -15216 9524
rect -15268 9452 -15216 9462
rect -14017 9512 -13965 9522
rect -16678 9440 -16626 9450
rect -16678 9378 -16626 9388
rect -16673 9086 -16630 9378
rect -16678 9076 -16626 9086
rect -16678 9014 -16626 9024
rect -17793 8550 -17792 8602
rect -17740 8550 -17739 8602
rect -17793 8548 -17739 8550
rect -17792 8530 -17740 8548
rect -19195 8238 -19143 8248
rect -19195 8176 -19143 8186
rect -20340 7803 -20288 7813
rect -20340 7741 -20288 7751
rect -19767 7805 -19715 7815
rect -19192 7803 -19146 8176
rect -19715 7755 -19145 7803
rect -19767 7743 -19715 7753
rect -20335 7429 -20291 7741
rect -20339 7419 -20287 7429
rect -20339 7357 -20287 7367
rect -21155 6981 -21102 6991
rect -21155 6917 -21102 6927
rect -20446 6989 -20393 6999
rect -20446 6925 -20393 6935
rect -21152 6433 -21106 6917
rect -21157 6423 -21102 6433
rect -21157 6358 -21102 6368
rect -20441 6140 -20397 6925
rect -20361 6875 -20308 6885
rect -20361 6811 -20308 6821
rect -20357 6226 -20313 6811
rect -19205 6594 -19152 6604
rect -19205 6530 -19152 6540
rect -20362 6216 -20309 6226
rect -19201 6224 -19156 6530
rect -20362 6151 -20309 6161
rect -19206 6214 -19153 6224
rect -20447 6130 -20393 6140
rect -20447 6064 -20393 6074
rect -20357 5929 -20313 6151
rect -19206 6150 -19153 6160
rect -16674 6157 -16631 9014
rect -16526 8977 -16483 9450
rect -16531 8967 -16479 8977
rect -15262 8971 -15219 9452
rect -14017 9450 -13965 9460
rect -12566 9511 -12514 9521
rect -14011 8971 -13968 9450
rect -12566 9449 -12514 9459
rect -12762 9422 -12710 9432
rect -12762 9360 -12710 9370
rect -12758 9138 -12713 9360
rect -12762 9128 -12709 9138
rect -12762 9064 -12709 9074
rect -16531 8905 -16479 8915
rect -15268 8961 -15216 8971
rect -15268 8899 -15216 8909
rect -14016 8961 -13964 8971
rect -12561 8970 -12518 9449
rect -11314 9429 -11262 9439
rect -11314 9367 -11262 9377
rect -14016 8899 -13964 8909
rect -12567 8960 -12515 8970
rect -12567 8898 -12515 8908
rect -11309 8804 -11266 9367
rect -11314 8794 -11262 8804
rect -11314 8732 -11262 8742
rect -15303 6872 -15251 6882
rect -15303 6810 -15251 6820
rect -15300 6449 -15254 6810
rect -16679 6147 -16626 6157
rect -16679 6083 -16626 6093
rect -20361 5919 -20308 5929
rect -20361 5854 -20308 5864
rect -19789 4561 -19736 4571
rect -19789 4496 -19736 4506
rect -19867 3896 -19822 3908
rect -19871 3886 -19818 3896
rect -19871 3821 -19818 3831
rect -19785 3823 -19740 4496
rect -15299 4204 -15255 6449
rect -16668 4185 -16614 4195
rect -17339 4153 -17286 4163
rect -16668 4119 -16614 4129
rect -15987 4191 -15933 4201
rect -15987 4126 -15933 4136
rect -15304 4194 -15250 4204
rect -15304 4128 -15250 4138
rect -17339 4088 -17286 4098
rect -19864 3567 -19828 3821
rect -19873 3557 -19820 3567
rect -19873 3492 -19820 3502
rect -17337 3469 -17288 4088
rect -17339 3459 -17286 3469
rect -16664 3466 -16615 4119
rect -15985 3469 -15935 4126
rect -17339 3393 -17286 3403
rect -16666 3456 -16612 3466
rect -15985 3463 -15931 3469
rect -15301 3468 -15251 4128
rect -16666 3390 -16612 3400
rect -15984 3459 -15931 3463
rect -15984 3394 -15931 3404
rect -15304 3458 -15251 3468
rect -15304 3393 -15251 3403
use sky130_fd_pr__nfet_01v8_lvt_93KYW7  XM1
timestamp 1659038648
transform 0 -1 -20745 1 0 5149
box -896 -310 896 310
use sky130_fd_pr__nfet_01v8_lvt_93KYW7  XM2
timestamp 1659038648
transform 0 -1 -20099 1 0 5149
box -896 -310 896 310
use sky130_fd_pr__pfet_01v8_lvt_PENQFR  XM3
timestamp 1659038648
transform 1 0 -18467 0 1 8028
box -496 -1337 496 1337
use sky130_fd_pr__pfet_01v8_lvt_PENQFR  XM4
timestamp 1659038648
transform 1 0 -14710 0 1 8028
box -496 -1337 496 1337
use sky130_fd_pr__pfet_01v8_lvt_UQCWFZ  XM5
timestamp 1659038648
transform 1 0 -13362 0 1 8028
box -596 -1337 596 1337
use sky130_fd_pr__pfet_01v8_lvt_CENSV5  XM6
timestamp 1659038648
transform 1 0 -19713 0 1 6954
box -496 -719 496 719
use sky130_fd_pr__nfet_01v8_lvt_L9TQ3V  XM7
timestamp 1659110821
transform 1 0 -18240 0 1 4763
box -296 -1319 296 1319
use sky130_fd_pr__nfet_01v8_lvt_L9TQ3V  XM8
timestamp 1659110821
transform 1 0 -16966 0 1 4763
box -296 -1319 296 1319
use sky130_fd_pr__pfet_01v8_lvt_5V5YF9  XM9
timestamp 1659038648
transform -1 0 -20759 0 -1 8028
box -296 -1337 296 1337
use sky130_fd_pr__pfet_01v8_lvt_PENQFR  XM10
timestamp 1659038648
transform 1 0 -17202 0 1 8028
box -496 -1337 496 1337
use sky130_fd_pr__nfet_01v8_lvt_L9TQ3V  XM11
timestamp 1659110821
transform 1 0 -19424 0 1 4763
box -296 -1319 296 1319
use sky130_fd_pr__pfet_01v8_lvt_PENQFR  XM12
timestamp 1659038648
transform 1 0 -15956 0 1 8028
box -496 -1337 496 1337
use sky130_fd_pr__pfet_01v8_lvt_UQCWFZ  XM14
timestamp 1659038648
transform 1 0 -11916 0 1 8028
box -596 -1337 596 1337
use sky130_fd_pr__pfet_01v8_lvt_CENSV5  XM19
timestamp 1659038648
transform 1 0 -19713 0 1 8646
box -496 -719 496 719
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ1 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1644243811
transform 1 0 -20690 0 1 3456
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ2
timestamp 1644243811
transform 1 0 -14620 0 1 3921
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ3
timestamp 1644243811
transform 1 0 -13822 0 1 3921
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ4
timestamp 1644243811
transform 1 0 -13024 0 1 3921
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ5
timestamp 1644243811
transform 1 0 -12226 0 1 3921
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ6
timestamp 1644243811
transform 1 0 -14628 0 1 3123
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ7
timestamp 1644243811
transform 1 0 -13830 0 1 3123
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ8
timestamp 1644243811
transform 1 0 -13032 0 1 3123
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ9
timestamp 1644243811
transform 1 0 -12234 0 1 3123
box 0 0 796 796
use sky130_fd_pr__res_xhigh_po_1p41_BPA34M  XR1
timestamp 1659038648
transform 0 -1 -13207 1 0 6231
box -307 -1378 307 1378
use sky130_fd_pr__res_xhigh_po_1p41_BPA34M  XR2
timestamp 1659038648
transform 1 0 -20748 0 1 2084
box -307 -1378 307 1378
use sky130_fd_pr__res_xhigh_po_1p41_BPA34M  XR3
timestamp 1659038648
transform -1 0 -20152 0 -1 2084
box -307 -1378 307 1378
use sky130_fd_pr__res_xhigh_po_1p41_BPA34M  XR4
timestamp 1659038648
transform 1 0 -19538 0 1 2084
box -307 -1378 307 1378
use sky130_fd_pr__res_xhigh_po_1p41_BPA34M  XR5
timestamp 1659038648
transform -1 0 -18942 0 -1 2084
box -307 -1378 307 1378
use sky130_fd_pr__res_xhigh_po_1p41_BPA34M  XR6
timestamp 1659038648
transform -1 0 -18346 0 -1 2084
box -307 -1378 307 1378
use sky130_fd_pr__res_xhigh_po_1p41_BPA34M  XR7
timestamp 1659038648
transform -1 0 -17750 0 -1 2084
box -307 -1378 307 1378
use sky130_fd_pr__res_xhigh_po_1p41_BPA34M  XR8
timestamp 1659038648
transform -1 0 -17154 0 -1 2084
box -307 -1378 307 1378
use sky130_fd_pr__res_xhigh_po_1p41_BPA34M  XR9
timestamp 1659038648
transform -1 0 -16558 0 -1 2084
box -307 -1378 307 1378
use sky130_fd_pr__res_xhigh_po_1p41_BPA34M  XR10
timestamp 1659038648
transform -1 0 -15962 0 -1 2084
box -307 -1378 307 1378
use sky130_fd_pr__res_xhigh_po_1p41_BPA34M  XR11
timestamp 1659038648
transform -1 0 -15366 0 -1 2084
box -307 -1378 307 1378
use sky130_fd_pr__res_xhigh_po_1p41_BPA34M  XR12
timestamp 1659038648
transform 0 -1 -13699 1 0 2824
box -307 -1378 307 1378
use sky130_fd_pr__res_xhigh_po_1p41_BPA34M  XR13
timestamp 1659038648
transform 0 -1 -13698 1 0 2228
box -307 -1378 307 1378
use sky130_fd_pr__res_xhigh_po_1p41_BPA34M  XR14
timestamp 1659038648
transform 0 -1 -13699 1 0 1632
box -307 -1378 307 1378
use sky130_fd_pr__res_xhigh_po_1p41_BPA34M  XR15
timestamp 1659038648
transform 0 -1 -13699 1 0 1036
box -307 -1378 307 1378
use sky130_fd_pr__res_xhigh_po_1p41_BPA34M  XR16
timestamp 1659038648
transform 1 0 -12031 0 1 1753
box -307 -1378 307 1378
use sky130_fd_pr__res_xhigh_po_1p41_BPA34M  XR17
timestamp 1659038648
transform 0 1 -13698 -1 0 439
box -307 -1378 307 1378
use sky130_fd_pr__res_xhigh_po_1p41_BPA34M  XR18
timestamp 1659038648
transform 0 -1 -16441 1 0 417
box -307 -1378 307 1378
use sky130_fd_pr__res_xhigh_po_1p41_BPA34M  XR19
timestamp 1659038648
transform 0 -1 -19179 1 0 417
box -307 -1378 307 1378
use sky130_fd_pr__res_xhigh_po_1p41_BPA34M  XR20
timestamp 1659038648
transform 0 -1 -13209 1 0 5631
box -307 -1378 307 1378
use sky130_fd_pr__res_xhigh_po_1p41_BPA34M  XR21
timestamp 1659038648
transform 0 1 -13209 -1 0 5017
box -307 -1378 307 1378
use sky130_fd_pr__nfet_01v8_lvt_L9TQ3V  sky130_fd_pr__nfet_01v8_lvt_L9TQ3V_0
timestamp 1659110821
transform 1 0 -18832 0 1 4763
box -296 -1319 296 1319
use sky130_fd_pr__nfet_01v8_lvt_L9TQ3V  sky130_fd_pr__nfet_01v8_lvt_L9TQ3V_1
timestamp 1659110821
transform 1 0 -17648 0 1 4763
box -296 -1319 296 1319
use sky130_fd_pr__nfet_01v8_lvt_L9TQ3V  sky130_fd_pr__nfet_01v8_lvt_L9TQ3V_2
timestamp 1659110821
transform 1 0 -16292 0 1 4764
box -296 -1319 296 1319
use sky130_fd_pr__nfet_01v8_lvt_L9TQ3V  sky130_fd_pr__nfet_01v8_lvt_L9TQ3V_3
timestamp 1659110821
transform 1 0 -15614 0 1 4764
box -296 -1319 296 1319
use sky130_fd_pr__nfet_01v8_lvt_L9TQ3V  sky130_fd_pr__nfet_01v8_lvt_L9TQ3V_4
timestamp 1659110821
transform 1 0 -14916 0 1 4764
box -296 -1319 296 1319
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VREF
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 VDD
port 2 nsew
<< end >>
