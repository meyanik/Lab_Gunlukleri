magic
tech sky130A
magscale 1 2
timestamp 1659038648
<< nwell >>
rect -296 -1337 296 1337
<< pmoslvt >>
rect -100 118 100 1118
rect -100 -1118 100 -118
<< pdiff >>
rect -158 1106 -100 1118
rect -158 130 -146 1106
rect -112 130 -100 1106
rect -158 118 -100 130
rect 100 1106 158 1118
rect 100 130 112 1106
rect 146 130 158 1106
rect 100 118 158 130
rect -158 -130 -100 -118
rect -158 -1106 -146 -130
rect -112 -1106 -100 -130
rect -158 -1118 -100 -1106
rect 100 -130 158 -118
rect 100 -1106 112 -130
rect 146 -1106 158 -130
rect 100 -1118 158 -1106
<< pdiffc >>
rect -146 130 -112 1106
rect 112 130 146 1106
rect -146 -1106 -112 -130
rect 112 -1106 146 -130
<< nsubdiff >>
rect -260 1267 -164 1301
rect 164 1267 260 1301
rect -260 1205 -226 1267
rect 226 1205 260 1267
rect -260 -1267 -226 -1205
rect 226 -1267 260 -1205
rect -260 -1301 -164 -1267
rect 164 -1301 260 -1267
<< nsubdiffcont >>
rect -164 1267 164 1301
rect -260 -1205 -226 1205
rect 226 -1205 260 1205
rect -164 -1301 164 -1267
<< poly >>
rect -100 1199 100 1215
rect -100 1165 -84 1199
rect 84 1165 100 1199
rect -100 1118 100 1165
rect -100 71 100 118
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -118 100 -71
rect -100 -1165 100 -1118
rect -100 -1199 -84 -1165
rect 84 -1199 100 -1165
rect -100 -1215 100 -1199
<< polycont >>
rect -84 1165 84 1199
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -1199 84 -1165
<< locali >>
rect -260 1267 -164 1301
rect 164 1267 260 1301
rect -260 1205 -226 1267
rect 226 1205 260 1267
rect -100 1165 -84 1199
rect 84 1165 100 1199
rect -146 1106 -112 1122
rect -146 114 -112 130
rect 112 1106 146 1122
rect 112 114 146 130
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -130 -112 -114
rect -146 -1122 -112 -1106
rect 112 -130 146 -114
rect 112 -1122 146 -1106
rect -100 -1199 -84 -1165
rect 84 -1199 100 -1165
rect -260 -1267 -226 -1205
rect 226 -1267 260 -1205
rect -260 -1301 -164 -1267
rect 164 -1301 260 -1267
<< viali >>
rect -84 1165 84 1199
rect -146 130 -112 1106
rect 112 130 146 1106
rect -84 37 84 71
rect -84 -71 84 -37
rect -146 -1106 -112 -130
rect 112 -1106 146 -130
rect -84 -1199 84 -1165
<< metal1 >>
rect -96 1199 96 1205
rect -96 1165 -84 1199
rect 84 1165 96 1199
rect -96 1159 96 1165
rect -152 1106 -106 1118
rect -152 130 -146 1106
rect -112 130 -106 1106
rect -152 118 -106 130
rect 106 1106 152 1118
rect 106 130 112 1106
rect 146 130 152 1106
rect 106 118 152 130
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect -152 -130 -106 -118
rect -152 -1106 -146 -130
rect -112 -1106 -106 -130
rect -152 -1118 -106 -1106
rect 106 -130 152 -118
rect 106 -1106 112 -130
rect 146 -1106 152 -130
rect 106 -1118 152 -1106
rect -96 -1165 96 -1159
rect -96 -1199 -84 -1165
rect 84 -1199 96 -1165
rect -96 -1205 96 -1199
<< properties >>
string FIXED_BBOX -243 -1284 243 1284
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 5.0 l 1.0 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
