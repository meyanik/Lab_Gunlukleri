magic
tech sky130A
magscale 1 2
timestamp 1659001593
<< nwell >>
rect 1584 1218 1643 1229
rect 1583 1161 1643 1218
rect 1583 1153 1642 1161
rect 1611 1135 1612 1153
rect 1597 923 1612 1135
rect 1597 884 1630 923
<< pwell >>
rect 1693 233 1702 263
rect 680 61 973 146
rect 2020 62 2121 391
rect 737 -252 765 61
rect 1761 27 2121 62
rect 1142 -26 1259 -24
rect 1142 -27 1193 -26
rect 1142 -75 1170 -27
rect 1229 -75 1259 -26
rect 1465 -48 1639 -37
rect 1465 -63 1674 -48
rect 1500 -84 1674 -63
rect 737 -314 1106 -252
rect 2020 -383 2121 27
rect 1281 -434 2146 -383
rect 1281 -436 1951 -434
rect 2020 -436 2121 -434
<< viali >>
rect 826 951 864 1191
rect 1143 1118 1177 1321
rect 1507 1124 1541 1327
rect 845 -78 879 264
rect 1160 132 1195 280
rect 1551 195 1585 277
<< metal1 >>
rect 680 1747 1393 1749
rect 680 1746 1436 1747
rect 680 1693 1397 1746
rect 1450 1693 1460 1746
rect 681 1691 1436 1693
rect 404 1111 604 1223
rect 681 1111 746 1691
rect 1217 1575 1227 1628
rect 1280 1627 1290 1628
rect 1280 1626 1698 1627
rect 2066 1626 2096 1628
rect 1280 1575 2096 1626
rect 1677 1574 2096 1575
rect 966 1389 1714 1460
rect 1137 1321 1183 1333
rect 1048 1213 1095 1239
rect 820 1191 870 1203
rect 904 1193 969 1196
rect 1048 1195 1105 1213
rect 820 1112 826 1191
rect 790 1111 826 1112
rect 404 1051 826 1111
rect 404 1023 604 1051
rect 790 1049 826 1051
rect 820 951 826 1049
rect 864 1112 870 1191
rect 903 1166 969 1193
rect 903 1112 938 1166
rect 1053 1159 1105 1195
rect 1058 1145 1105 1159
rect 864 1049 938 1112
rect 864 951 870 1049
rect 820 939 870 951
rect 903 905 938 1049
rect 970 940 1034 1110
rect 1074 1029 1105 1145
rect 1137 1118 1143 1321
rect 1177 1215 1183 1321
rect 1501 1327 1547 1339
rect 1501 1215 1507 1327
rect 1177 1181 1507 1215
rect 1177 1118 1183 1181
rect 1137 1106 1183 1118
rect 1501 1124 1507 1181
rect 1541 1124 1547 1327
rect 2066 1298 2096 1574
rect 1584 1218 1643 1229
rect 1583 1161 1643 1218
rect 1728 1205 2096 1298
rect 1583 1153 1642 1161
rect 1501 1112 1547 1124
rect 1074 1027 1290 1029
rect 1074 981 1229 1027
rect 1074 922 1105 981
rect 1219 975 1229 981
rect 1281 975 1291 1027
rect 903 863 963 905
rect 1057 883 1105 922
rect 1584 923 1612 1153
rect 1650 952 1719 1120
rect 916 861 963 863
rect 1052 852 1105 883
rect 1389 866 1399 918
rect 1451 914 1461 918
rect 1584 914 1630 923
rect 1451 904 1630 914
rect 1451 872 1653 904
rect 1451 866 1461 872
rect 1584 871 1653 872
rect 2066 851 2096 1205
rect 1723 758 2096 851
rect 1446 674 1720 681
rect 968 616 1720 674
rect 541 477 741 532
rect 1263 488 1335 616
rect 1446 612 1720 616
rect 2066 489 2096 758
rect 1216 477 1335 488
rect 541 465 1335 477
rect 1615 468 1738 469
rect 1615 465 1768 468
rect 541 413 1768 465
rect 541 332 741 413
rect 839 264 885 276
rect 494 146 694 208
rect 839 146 845 264
rect 494 61 845 146
rect 494 8 694 61
rect 737 -252 765 61
rect 839 -78 845 61
rect 879 146 885 264
rect 983 230 1060 413
rect 1216 412 1768 413
rect 1216 340 1288 412
rect 1645 411 1768 412
rect 1154 280 1201 292
rect 879 61 973 146
rect 1154 132 1160 280
rect 1195 264 1201 280
rect 1545 277 1591 289
rect 1545 264 1551 277
rect 1195 209 1551 264
rect 1195 132 1201 209
rect 1545 195 1551 209
rect 1585 195 1591 277
rect 1689 263 1765 411
rect 1941 289 2141 489
rect 1689 237 1803 263
rect 1693 233 1803 237
rect 1545 183 1591 195
rect 1154 120 1201 132
rect 1329 62 1339 119
rect 1408 118 1418 119
rect 1486 118 1589 119
rect 1634 118 1690 119
rect 1408 113 1690 118
rect 1408 86 1700 113
rect 1408 62 1696 86
rect 1444 61 1696 62
rect 879 -78 885 61
rect 1698 57 1700 86
rect 2020 62 2121 289
rect 1222 49 1232 57
rect 1047 11 1232 49
rect 1222 4 1232 11
rect 1285 48 1295 57
rect 1285 12 1300 48
rect 1761 27 2121 62
rect 1285 4 1295 12
rect 1142 -28 1312 -24
rect 839 -90 885 -78
rect 987 -37 1380 -28
rect 1699 -37 1760 -31
rect 987 -87 1760 -37
rect 987 -88 1473 -87
rect 1154 -89 1201 -88
rect 952 -252 1334 -251
rect 737 -313 1334 -252
rect 1408 -313 1419 -251
rect 737 -314 1106 -313
rect 2020 -383 2121 27
rect 1281 -384 2146 -383
rect 1220 -436 1230 -384
rect 1285 -434 2146 -384
rect 1285 -436 1951 -434
rect 2020 -436 2121 -434
<< via1 >>
rect 1397 1693 1450 1746
rect 1227 1575 1280 1628
rect 1229 975 1281 1027
rect 1399 866 1451 918
rect 1339 62 1408 119
rect 1232 4 1285 57
rect 1334 -313 1408 -251
rect 1230 -436 1285 -384
<< metal2 >>
rect 1397 1746 1450 1756
rect 1397 1683 1450 1693
rect 1227 1628 1280 1638
rect 1227 1565 1280 1575
rect 1228 1037 1280 1565
rect 1399 1564 1448 1683
rect 1228 1027 1281 1037
rect 1228 982 1229 1027
rect 1229 965 1281 975
rect 1399 918 1451 1564
rect 1399 856 1451 866
rect 1339 123 1408 129
rect 1333 119 1411 123
rect 1232 63 1285 67
rect 1231 57 1286 63
rect 1231 4 1232 57
rect 1285 4 1286 57
rect 1231 -356 1286 4
rect 1333 62 1339 119
rect 1408 62 1411 119
rect 1333 -6 1411 62
rect 1333 -37 1409 -6
rect 1333 -251 1411 -37
rect 1333 -294 1334 -251
rect 1408 -294 1411 -251
rect 1334 -323 1408 -313
rect 1230 -384 1286 -356
rect 1285 -404 1286 -384
rect 1230 -446 1285 -436
use sky130_fd_pr__nfet_01v8_648S5X  XM1
timestamp 1659001593
transform 1 0 1019 0 1 100
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  sky130_fd_pr__nfet_01v8_648S5X_0
timestamp 1659001593
transform 1 0 1726 0 1 100
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_UGSVTG  sky130_fd_pr__pfet_01v8_UGSVTG_0
timestamp 1659001593
transform 1 0 1003 0 1 1029
box -211 -537 211 537
use sky130_fd_pr__pfet_01v8_UGSVTG  sky130_fd_pr__pfet_01v8_UGSVTG_1
timestamp 1659001593
transform 1 0 1682 0 1 1040
box -211 -537 211 537
<< labels >>
flabel metal1 541 332 741 532 0 FreeSans 256 0 0 0 A
port 0 nsew
flabel metal1 404 1023 604 1223 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 1941 289 2141 489 0 FreeSans 256 0 0 0 O
port 2 nsew
flabel metal1 494 8 694 208 0 FreeSans 256 0 0 0 VSS
port 3 nsew
<< end >>
