** sch_path: /home/ubuntu/Desktop/design/xschem/inv_TB.sch
**.subckt inv_TB
X1 in VDD out GND inv
V1 in GND pulse 0 1.8 2n 1n 1n 10n 20n
V2 VDD GND 1.8
**** begin user architecture code

** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt_mm




.include ../netgen/inv_pex.spice
.control

save all

tran 0.1n 200n
write inv_TB.raw
plot v(out) v(in)+3
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
