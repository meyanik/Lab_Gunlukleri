magic
tech sky130A
magscale 1 2
timestamp 1659038648
<< nwell >>
rect -496 -1337 496 1337
<< pmoslvt >>
rect -300 118 300 1118
rect -300 -1118 300 -118
<< pdiff >>
rect -358 1106 -300 1118
rect -358 130 -346 1106
rect -312 130 -300 1106
rect -358 118 -300 130
rect 300 1106 358 1118
rect 300 130 312 1106
rect 346 130 358 1106
rect 300 118 358 130
rect -358 -130 -300 -118
rect -358 -1106 -346 -130
rect -312 -1106 -300 -130
rect -358 -1118 -300 -1106
rect 300 -130 358 -118
rect 300 -1106 312 -130
rect 346 -1106 358 -130
rect 300 -1118 358 -1106
<< pdiffc >>
rect -346 130 -312 1106
rect 312 130 346 1106
rect -346 -1106 -312 -130
rect 312 -1106 346 -130
<< nsubdiff >>
rect -460 1267 -364 1301
rect 364 1267 460 1301
rect -460 1205 -426 1267
rect 426 1205 460 1267
rect -460 -1267 -426 -1205
rect 426 -1267 460 -1205
rect -460 -1301 -364 -1267
rect 364 -1301 460 -1267
<< nsubdiffcont >>
rect -364 1267 364 1301
rect -460 -1205 -426 1205
rect 426 -1205 460 1205
rect -364 -1301 364 -1267
<< poly >>
rect -300 1199 300 1215
rect -300 1165 -284 1199
rect 284 1165 300 1199
rect -300 1118 300 1165
rect -300 71 300 118
rect -300 37 -284 71
rect 284 37 300 71
rect -300 21 300 37
rect -300 -37 300 -21
rect -300 -71 -284 -37
rect 284 -71 300 -37
rect -300 -118 300 -71
rect -300 -1165 300 -1118
rect -300 -1199 -284 -1165
rect 284 -1199 300 -1165
rect -300 -1215 300 -1199
<< polycont >>
rect -284 1165 284 1199
rect -284 37 284 71
rect -284 -71 284 -37
rect -284 -1199 284 -1165
<< locali >>
rect -460 1267 -364 1301
rect 364 1267 460 1301
rect -460 1205 -426 1267
rect 426 1205 460 1267
rect -300 1165 -284 1199
rect 284 1165 300 1199
rect -346 1106 -312 1122
rect -346 114 -312 130
rect 312 1106 346 1122
rect 312 114 346 130
rect -300 37 -284 71
rect 284 37 300 71
rect -300 -71 -284 -37
rect 284 -71 300 -37
rect -346 -130 -312 -114
rect -346 -1122 -312 -1106
rect 312 -130 346 -114
rect 312 -1122 346 -1106
rect -300 -1199 -284 -1165
rect 284 -1199 300 -1165
rect -460 -1267 -426 -1205
rect 426 -1267 460 -1205
rect -460 -1301 -364 -1267
rect 364 -1301 460 -1267
<< viali >>
rect -284 1165 284 1199
rect -346 130 -312 1106
rect 312 130 346 1106
rect -284 37 284 71
rect -284 -71 284 -37
rect -346 -1106 -312 -130
rect 312 -1106 346 -130
rect -284 -1199 284 -1165
<< metal1 >>
rect -296 1199 296 1205
rect -296 1165 -284 1199
rect 284 1165 296 1199
rect -296 1159 296 1165
rect -352 1106 -306 1118
rect -352 130 -346 1106
rect -312 130 -306 1106
rect -352 118 -306 130
rect 306 1106 352 1118
rect 306 130 312 1106
rect 346 130 352 1106
rect 306 118 352 130
rect -296 71 296 77
rect -296 37 -284 71
rect 284 37 296 71
rect -296 31 296 37
rect -296 -37 296 -31
rect -296 -71 -284 -37
rect 284 -71 296 -37
rect -296 -77 296 -71
rect -352 -130 -306 -118
rect -352 -1106 -346 -130
rect -312 -1106 -306 -130
rect -352 -1118 -306 -1106
rect 306 -130 352 -118
rect 306 -1106 312 -130
rect 346 -1106 352 -130
rect 306 -1118 352 -1106
rect -296 -1165 296 -1159
rect -296 -1199 -284 -1165
rect 284 -1199 296 -1165
rect -296 -1205 296 -1199
<< properties >>
string FIXED_BBOX -443 -1284 443 1284
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 5.0 l 3.0 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
